module mux_unstriping ();
endmodule